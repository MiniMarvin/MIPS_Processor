module mul (
	input clk,       // Clock
	input clk_en,    // Clock Enable
	input rst_n,     // Asynchronous reset active low
	input module_en, // Enable the operation of the module
	input start_div, // Start the 
	output ready,    // Inform that no division is occurring
	output quotient, // Quotient of the division
	output rest      // Rest of the division value
	
);

endmodule