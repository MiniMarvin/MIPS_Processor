module partControl (
	input clk,    // Clock
	input clk_en, // Clock Enable
	input rst_n,  // Asynchronous reset active low
	input ignore_amt   // Defines the amount of numbers to ignore
);

// Control wich part of the word is going to pass the other part is going to become zero


endmodule