module divMul (
	input clk,    // Clock
	input clk_en, // Clock Enable
	input rst_n,  // Asynchronous reset active low
	input divMul,  // Asynchronous reset active low
	output ready,
	output reg hi,
	output reg lo
);


// The magic box to div/mul



endmodule
